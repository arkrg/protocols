package apb_pkg;
    parameter int NUM_SLAVE = 4;
    parameter int ADDR_WIDTH = 12;
    parameter int DATA_WIDTH = 32;
endpackage
